// contant value memory
module M0
  (
   input [7:0] M0VAL,
   output [7:0] RDATA
   );
   assign RDATA = M0VAL;
   
endmodule // M0


